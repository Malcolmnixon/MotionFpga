--! @mainpage MachX02-7000HE MotionFPGA
--!
--! @section Introduction
--! This documentation describes the MotionFPGA for the MachX02-7000HE target.
--!
--! @section sec_top Top Component
--! Todo
--! @sa top

